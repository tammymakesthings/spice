Band-Pass Filter

Vin 1 0 DC 0 AC 1
C1 1 2 0.0001m
L1 2 3 1
R1 3 0 100

.AC LIN 1000 0.1 1000
.TRAN 	5US  500US
* VIEW RESULTS
.PRINT	AC 	VM(2) VP(2)
.PLOT	AC	VM(2) VP(2)
.PRINT	TRAN 	V(1) V(2)
.PLOT	TRAN 	V(1) V(2)
.PROBE
.end
